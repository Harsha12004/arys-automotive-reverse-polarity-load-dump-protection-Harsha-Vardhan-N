* Step 1: Basic NGspice Test Circuit

Vin in 0 DC 12
Rload in 0 100

.tran 1ms 20ms
.end

