* STEP 2 - Reverse Polarity Protection using Diode

Vin in 0 DC 12

* Reverse polarity protection diode
D1 in out Dmodel

.model Dmodel D(BV=40 IBV=1mA RS=0.1 TT=1u)

* Load
Rload out 0 100

.tran 1ms 40ms
.end
