* STEP 3 - Load Dump Protection with TVS Diode (Corrected)

Vin in 0 PWL(0 12  1m 12  2m 80  352m 80  353m 12)

* Reverse polarity diode (correct orientation)
D1 mid in Dmodel
.model Dmodel D(BV=40 IBV=1mA RS=0.1 TT=1u)

* TVS diode to clamp surge
D2 mid 0 TVS48
.model TVS48 D(BV=48 IBV=1m RS=0.05 CJO=200p)

* Load
Rload mid 0 100

.tran 0.1m 400m
.end
